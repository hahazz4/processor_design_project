module pc_increment();



endmodule