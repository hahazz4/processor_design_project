//Start of code

//Carry Look Ahead Adder
module carry_out(input reg [15:0] 
                  output [31:0] );
    
    always @(negedge clk){
        begin

        end
    }    
endmodule
//End of code