module shift_left_()

endmodule