module datapath();
    reg s;
    encoder ecode(s);
    multiplexer mplex(s);
endmodule //Register end.