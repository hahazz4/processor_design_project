module select_encode();