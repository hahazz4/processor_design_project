module rotate_right(input [31:0] A, r_num,
                           output [31:0] rotateR_result);

endmodule