`timescale 1ns/10ps
module control_unit(
    input [31:0] instruction_reg,
    input clk, reset, stop, …, con_ff,
    output reg Gra, Grb, Grc, R_enable, …, R_select, // define the inputs and outputs to your Control Unit
    Y_enable, Z_enable, PC_select, PC_increment_enable, …, MAR_enable,
    read, write, …, clr,
    ADD, AND, …, SHR,);

parameter Reset_state= 8'b00000000, fetch0 = 8'b00000001, fetch1 = 8'b00000010, fetch2= 8'b00000011,
          add3 = 8'b00000100, add4= 8'b00000101, add5= 8'b00000110, sub3 = 8'b00000111, sub4 = 8'b00001000, sub5 = 8'b00001001,
          mul3 = 8'b00001010, mul4 = 8'b00001011, mul5 = 8'b00001100, mul6 = 8'b00001101, div3 = 8'b00001110, div4 = 8'b00001111,
          div5 = 8'b00010000, div6 = 8'b00010001, or3 = 8'b00010010, or4 = 8'b00010011, or5 = 8'b00010100, and3 = 8'b00010101, 
          and4 = 8'b00010110, and5 = 8'b00010111, shl3 = 8'b00011000, shl4 = 8'b00011001, shl5 = 8'b00011010, shr3 = 8'b00011011,
          shr4 = 8'b00011100, shr5 = 8'b00011101, rol3 = 8'b00011110, rol4 = 8'b00011111, rol5 = 8'b00100000, ror3 = 8'b00100001,
          ror4 = 8'b00100010, ror5 = 8'b00100011, neg3 = 8'b00100100, neg4 = 8'b00100101, neg5 = 8'b00100110, not3 = 8'b00100111,
          not4 = 8'b00101000, not5 = 8'b00101001, ld3 = 8'b00101010, ld4 = 8'b00101011, ld5 = 8'b00101100, ld6 = 8'b00101101, 
          ld7 = 8'b00101110, ldi3 = 8'b00101111, ldi4 = 8'b00110000, ldi5 = 8'b00110001, st3 = 8'b00110010, st4 = 8'b00110011,
          st5 = 8'b00110100, st6 = 8'b00110101, st7 = 8'b00110110, addi3 = 8'b00110111, addi4 = 8'b00111000, addi5 = 8'b00111001,
          andi3 = 8'b00111010, andi4 = 8'b00111011, andi5 = 8'b00111100, ori3 = 8'b00111101, ori4 = 8'b00111110, ori5 = 8'b00111111,
          br3 = 8'b01000000, br4 = 8'b01000001, br5 = 8'b01000010, br6 = 8'b01000011, br7 = 8'b11111111, jr3 = 8'b01000100, jal3 = 8'b01000101, 
          jal4 = 8'b01000110, mfhi3 = 8'b01000111, mflo3 = 8'b01001000, in3 = 8'b01001001, out3 = 8'b01001010, nop3 = 8'b01001011, 
          halt3 = 8'b01001100;

//    addition_op = 5'b00011, 
//    subtraction_op = 5'b00100, 
//    multiplication_op = 5'b01111, 
//    division_op = 5'b10000, 
//    left_shift_op = 5'b01001, 
//    right_shift_op = 5'b00111, 
//    arith_shift_right_op = 5'b01000, 
//    left_rotate_op = 5'b01011, 
//    right_rotate_op = 5'b01010, 
//    and_op = 5'b00101, 
//    or_op = 5'b00110, 
//    negate_op = 5'b10001, 
//    not_op = 5'b10010;
//    ldw_op = 5'b00000;
//    ldi_op = 5'b00001;
//    stw_op = 5'b00010;
//    addi_op = 5'b01100;
//    andi_op = 5'b01100;
//    ori_op = 5'b01110;
//    br_op = 5'b10011;
//    // brzr_op = 5'b10011;
//    // brnz_op = 5'b10011;
//    // brmi_op = 5'b10011;
//    // brpl_op = 5'b10011;
//    jr_op = 5'b10100;
//    jal_op = 5'b10101;
//    mfhi_op = 5'b11000;
//    mflo_op = 5'b11001;
//    out = 5'b10111;
//    in = 5'b10110;
//    nop = 5'b11010;
//    halt = 5'b11011;

reg [7:0] present_state = reset_state;      // adjust the bit pattern based on the number of states

always @(posedge clk, posedge reset, posedge stop)  //con_ff finite state machine; if clk or reset rising-edge
begin
    if (Reset == 1'b1) present_state = reset_state;
    else case (present_state)
        reset_state : present_state = fetch0;
        fetch0 : present_state = fetch1;
        fetch1 : present_state = fetch2;
        fetch2 : begin
        case (instruction_reg [31:27]) // inst. decoding based on the opcode to set the next state
            5'b00011 : present_state = add3; 
            5'b00100 : present_state = sub3;
            5'b01111 : present_state = mul3;
            5'b10000 : present_state = div3;
            5'b00111 : present_state = shr3;
            5'b01001 : present_state = shl3;
            5'b01010 : present_state = ror3;
            5'b01011 : present_state = rol3;
            5'b00101 : present_state = and3;
            5'b00110 : present_state = or3;
            5'b10001 : present_state = neg3;
            5'b10010 : present_state = not3;
            5'b00000 : present_state = ld3;
            5'b00001 : present_state = ldi3;
            5'b00010 : present_state = st3;
            5'b01100 : present_state = addi3;
            5'b01100 : present_state = andi3;
            5'b01110 : present_state = ori3;
            5'b10011 : present_state = br3;
            5'b10100 : present_state = jr3;
            5'b10101 : present_state = jal3;
            5'b11000 : present_state = mfhi3;
            5'b11001 : present_state = mflo3;
            5'b10110 : present_state = in3;
            5'b10111 : present_state = out3;                
            5'b11010 : present_state = nop3;
            5'b11011 : present_state = halt3;
        endcase
        end

        add3 : Present_state = add4;
        add4 : Present_state = add5;
        add5 : Present_state = fetch0;
                
        addi3 : Present_state = addi4;
        addi4 :	Present_state = addi5;
        addi5 : Present_state = fetch0;
                
        sub3 : Present_state = sub4;
        sub4 : Present_state = sub5;
        sub5 : Present_state = fetch0;
        
        mul3 : Present_state = mul4;
        mul4 : Present_state = mul5;
        mul5 : Present_state = mul6;
        mul6 : Present_state = fetch0; 
        
        div3 : Present_state = div4;
        div4 : Present_state = div5;
        div5 : Present_state = div6;
        div6 : Present_state = fetch0;
                
        or3 : Present_state = or4;
        or4 : Present_state = or5;
        or5	: Present_state = fetch0;
                
        and3 : Present_state = and4;
        and4 : Present_state = and5;
        and5 : Present_state = fetch0;
                
        shl3 : Present_state = shl4;
        shl4 : Present_state = shl5;
        shl5 : Present_state = fetch0;
                
        shr3 : Present_state = shr4;
        shr4 : Present_state = shr5;
        shr5 : Present_state = fetch0;
                
        rol3 : Present_state = rol4;
        rol4 : Present_state = rol5;
        rol5 : Present_state = fetch0;
                
        ror3 : Present_state = ror4;
        ror4 : Present_state = ror5;
        ror5 : Present_state = fetch0;
                
        neg3 : Present_state = neg4;
        neg4 : Present_state = fetch0;
                
        not3 : Present_state = not4;
        not4 : Present_state = fetch0;
                
        ld3 : Present_state = ld4;
        ld4 : Present_state = ld5;
        ld5 : Present_state = ld6;
        ld6 : Present_state = ld7;
        ld7 : Present_state = fetch0;
                
        ldi3 : Present_state = ldi4;
        ldi4 : Present_state = ldi5;
        ldi5 : Present_state = fetch0;
                
        st3 : Present_state = st4;
        st4 : Present_state = st5;
        st5 : Present_state = st6;
        st6 : Present_state = st7;
        st7 : Present_state = fetch0;
                
        andi3 : Present_state = andi4;
        andi4 : Present_state = andi5;
        andi5 : Present_state = fetch0;
                
        ori3 : Present_state = ori4;
        ori4 : Present_state = ori5;
        ori5 : Present_state = fetch0;
                
        jal3 : Present_state = jal4;
        jal4 : Present_state = fetch0;
                
        jr3 : Present_state = fetch0;
                
        br3 : Present_state = br4;
        br4 : Present_state = br5;
        br5 : Present_state = br6;
        br6 : Present_state = br7;
        br7 : Present_state = fetch0;
                
        out3 : Present_state = fetch0;
                
        in3 : Present_state = fetch0;
                
        mflo3 : Present_state = fetch0;
        
        mfhi3 : Present_state = fetch0;
        
        nop3 : Present_state = fetch0;
    endcase
end

always @(present_state) // do the job for each state
begin
    case (present_state) // assert the requinstruction_reged signals in each state
    reset_state: begin
        Gra <= 0; Grb <= 0; Grc <= 0; Y_enable <= 0; PC_select <= 0; ZHighout <= 0; ZLowout <= 0; MDR_select <= 0; 
        MAR_enable <= 0; PC_enable <= 0; MDR_enable <= 0; instruction_reg_enable <= 0; Y_enable <= 0; PC_increment_enable <= 0; MDR_read <= 0;
		HIin <= 0; LOin <= 0; HIout <= 0; LOout <= 0; ZHighIn <= 0; ZLowIn <= 0; Cout <= 0; RAM_write <= 0; R_enable <= 0;
        R_select <= 0; BAout <= 0; CON_enable <= 0; enableInputPort <= 0; OutPort_enable <= 0; InPortout <= 0;
    end
    
    fetch0: begin
        PC_select <= 1; // see if you need to de-assert these signals
        MAR_enable <= 1;
        PC_increment_enable <= 1;
        Z_enable <= 0;
    end

	fetch1: begin
		PC_select <= 0; MAR_enable <= 0; 
		MDR_enable <= 1; MDR_read <= 1; ZLowout <= 1;
	end

	fetch2: begin
		MDR_enable <= 0; MDR_read <= 0; ZLowout <= 0;
		MDR_select <= 1; instruction_reg_enable <= 1; PC_enable <= 1; PC_increment_enable <= 1;	
		#21 PC_enable <= 0;
	end 

	//Add, Subtraction Operations
	add3, sub3: begin	
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;
		Grb <= 1; R_select <= 1; Y_enable <= 1;
	end

	add4, sub4: begin
		Grb <= 0; R_select <= 0; Y_enable <= 0;
		Grc <= 1; R_select <= 1; ZHighIn <= 1; ZLowIn <= 1; 
	end

	add5, sub5: begin
		Grc <= 0; R_select <= 0; ZHighIn <= 0; ZLowIn <= 0;
		ZLowout <= 1; Gra <= 1; R_enable <= 1;
	end

	//Or, And, Shift-Left, Shift-Right, Rotate-Left, Rotate-Right Operations
	or3, and3, shl3, shr3, rol3, ror3: begin	
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;
		Grb <= 1; R_select <= 1; Y_enable <= 1;
	end
	
    or4, and4, shl4, shr4, rol4, ror4: begin
		Grb <= 0; R_select <= 0; Y_enable <= 0;
		Grc <= 1; R_select <= 1; ZHighIn <= 1; ZLowIn <= 1;
	end
	
    or5, and5, shl5, shr5, rol5, ror5: begin
		Grc <= 0; R_select <= 0; ZHighIn <= 0;  ZLowIn <= 0;
		ZLowout <= 1; Gra <= 1; R_enable <= 1;
		#40 ZLowout <= 0; Gra <= 1; R_select <= 1; R_enable <= 0;
	end
		
    //Multiplication, Division Operations
	mul3, div3: begin	
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;
		Grb <= 1; R_select <= 1; Y_enable <= 1;  		
	end
	
    mul4, div4: begin
		Grb <= 0; R_select <= 0; Y_enable <= 0;
		Grc <= 1; R_select <= 1; ZHighIn <= 1; ZLowIn <= 1;			
	end
	
    mul5, div5: begin
		Grb <= 0; R_select <= 0; ZHighIn <= 0; ZLowIn <= 0;
		ZLowout <= 1; LOin <= 1;			
	end
	
    mul6, div6: begin
		ZLowout <= 0; LOin <= 0;
		ZHighout <= 1; HIin <= 1;
	end
		
    //Not, Negate Operations
	not3, neg3: begin	
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;
		Grb <= 1; R_select <= 1; ZHighIn <= 1; ZLowIn <= 1;
	end
	
    not4, neg4: begin
		Grb <= 0; R_select <= 0; ZHighIn <= 0; ZLowIn <= 0;
		ZLowout <= 1; Gra <= 1; R_enable <= 1;
	end

	//And Immediate Operation
	andi3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;	
		Grb <= 1; R_select <= 1; Y_enable <= 1;
	end

	andi4: begin
		Grb <= 0; R_select <= 0; Y_enable <= 0;
		Cout <= 1; ZHighIn <= 1; ZLowIn <= 1;
	end

	andi5: begin
		Cout <= 0; ZHighIn <= 0; ZLowIn <= 0;
		ZLowout <= 1; Gra <= 1; R_enable <= 1;
		#40 ZLowout <= 0; Gra <= 1; R_select <= 1; R_enable <= 0;
	end
		
    //Add Immediate Operation
	addi3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;	
		Grb <= 1; R_select <= 1; Y_enable <= 1;
	end

	addi4: begin
		Grb <= 0; R_select <= 0; Y_enable <= 0;
		Cout <= 1; ZHighIn <= 1;  ZLowIn <= 1;
	end

	addi5: begin
		Cout <= 0; ZHighIn <= 0;  ZLowIn <= 0;
		ZLowout <= 1; Gra <= 1; R_enable <= 1;
		#40 ZLowout <= 0; Gra <= 1; R_select <= 1; R_enable <= 0;
	end
		
    //Or Immediate Operation
	ori3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;		
		Grb <= 1; R_select <= 1; Y_enable <= 1;
	end

	ori4: begin
		Grb <= 0; R_select <= 0; Y_enable <= 0;
		Cout <= 1; ZHighIn <= 1;  ZLowIn <= 1;
	end

	ori5: begin
		Cout <= 0; ZHighIn <= 0;  ZLowIn <= 0;
		ZLowout <= 1; Gra <=1 ; R_enable <= 1;
		#40 ZLowout <= 0; Gra <= 1; R_select <= 1; R_enable <= 0;
	end
		
    //Load Operation
	ld3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;	
		Grb <= 1; BAout <= 1; Y_enable <= 1;
	end

	ld4: begin
		Grb <= 0; BAout <= 0; Y_enable <= 0;
		Cout <= 1; ZHighIn <= 1; ZLowIn <= 1;
	end

	ld5: begin
		Cout <= 0; ZHighIn <= 0;  ZLowIn <= 0;
		ZLowout <= 1; MAR_enable <= 1;
	end

	ld6: begin
		ZLowout <= 0; MAR_enable <= 0;
		MDR_read <= 1; MDR_enable <= 1;
	end
	
    ld7: begin
		MDR_read <= 0; MDR_enable <= 0;
		MDR_select <= 1; Gra <= 1; R_enable <= 1;
	end
		
    //Load Immediate Operation
	ldi3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;			
		Grb <= 1; BAout <= 1; Y_enable <= 1;
	end

	ldi4: begin
		Grb <= 0; BAout <= 0; Y_enable <= 0;
		Cout <=1; ZHighIn <= 1; ZLowIn <= 1;
	end

	ldi5: begin
		Cout <= 0; ZHighIn <= 0; ZLowIn <= 0;
		ZLowout <= 1; Gra <= 1; R_enable <= 1;
		#40 ZLowout <= 0; Gra <= 0; R_enable <= 0; 
	end
		
    //Store Operation
	st3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;		
		Grb <= 1; BAout <= 1; Y_enable <= 1;
	end

	st4: begin
		Grb <= 0; BAout <= 0; Y_enable <= 0;
		Cout <= 1; ZHighIn <= 1; ZLowIn <= 1;
	end

	st5: begin
		Cout <= 0; ZHighIn <= 0; ZLowIn <= 0;
		ZLowout <= 1; MAR_enable <= 1;
	end

	st6: begin
		ZLowout <= 0; MAR_enable <= 0;
		MDR_read <= 0; Gra <= 1; R_select <= 1; MDR_enable <= 1;
	end
	
    st7: begin
		Gra <= 0; R_select <= 0; MDR_enable <= 0;
		MDR_select <= 1; 
		#5 RAM_write <= 1; 
	end
		
    //Jump Register Operation
	jr3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;				
		Gra <= 1; R_select <= 1; PC_enable <= 1;
		#40 PC_enable <= 0;
	end
		
    //Jump and Link Operation
	jal3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;	
		PC_select <= 1; R_enableIn <= 16'h4000; 
	end

	jal4: begin
		R_enableIn <= 16'h0000; PC_select <= 0;		
		Gra <= 1; R_select <= 1; PC_enable <= 1;
	end
		
    //Move from Hi Register Operation
	mfhi3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;	
		Gra <= 1; R_enable <= 1; HIout <= 1;
		#40 Gra <= 0; R_enable <= 0; HIout <= 0;
	end
		
    //Move from Lo Register Operation
	mflo3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;	
		Gra <= 1; R_enable <= 1; LOout <= 1;
		#40 Gra <= 0; R_enable <= 0; LOout <= 0;
	end
		
    //Inputting Operation
	in3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;
		Gra <= 1; R_enable <= 1; InPortout <= 1;
	end
		
    //Outputting Operation
	out3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;	
		Gra <= 1; R_select <= 1; Y_enable <= 1; OutPort_enable <= 1;
	end
		
    //Branch Operation
	br3: begin
		MDR_select <= 0; instruction_reg_enable <= 0; PC_enable <= 0; PC_increment_enable <= 0;		
		Gra <= 1; R_select <= 1; CON_enable <= 1;
	end

	br4: begin
		Gra <= 0; R_select <= 0; CON_enable <= 0;
		PC_select <= 1; Y_enable <= 1;
	end

	br5: begin
		PC_select <= 0; Y_enable <= 0;
	   	Cout <= 1; ZHighIn <= 1; ZLowIn <= 1;
	end

	br6: begin
		Cout <= 0; ZHighIn <= 0; ZLowIn <= 0;
	   	ZLowout <= 1; PC_enable <= 1;
	end
	
    br7: begin
		ZLowout <= 0; PC_enable <= 0;
		PC_select <= 1; 
	end
		
    //No Operation
	nop3: begin
	end
		
    //Halt Operation (Stops instruction execution)
	halt3: begin
		Run <= 0;
	end
		
    //Any other input would be default to do nothing
    default: begin 
	end
    endcase
end
endmodule
