module memory_datapath(input clk, input clr, input MAR_enable, input MDR_enable, input read, input write, );

endmodule