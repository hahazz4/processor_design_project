module rotate_left(input [31:0] A, r_num,
                           output [31:0] rotateL_result);

endmodule